----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:01:10 03/29/2014 
-- Design Name: 
-- Module Name:    elevatorlogic - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity elevatorlogic is
    Port ( SW0 : in  STD_LOGIC;
           SW1 : in  STD_LOGIC;
           EN : in  STD_LOGIC;
           OUT0 : out  STD_LOGIC;
           OUT1 : out  STD_LOGIC);
end elevatorlogic;

architecture Behavioral of elevatorlogic is

begin


end Behavioral;

